module interrupt_handler (
    
); 
    
endmodule