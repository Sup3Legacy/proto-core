`define i_ 